/* Copyright(C) 2016 Cobac.Net All Rights Reserved. */
/* chapter: ��9�͉ۑ�       */
/* project: display_XGA     */
/* outline: XGA�p�p�����[�^ */

/* XGA(1024�~768)�p�����[�^ */
//localparam HPERIOD = 11'd1344;
//localparam HFRONT  = 11'd24;
//localparam HWIDTH  = 11'd136;
//localparam HBACK   = 11'd160;

//localparam VPERIOD = 10'd806;
//localparam VFRONT  = 10'd3;
//localparam VWIDTH  = 10'd6;
//localparam VBACK   = 10'd29;

/* FHD(1920*1080)�p�����[�^*/
localparam HPERIOD = 12'd2080;
localparam HFRONT  = 12'd48;
localparam HWIDTH  = 12'd32;
localparam HBACK   = 12'd80;

localparam VPERIOD = 11'd1111;
localparam VFRONT  = 11'd3;
localparam VWIDTH  = 11'd5;
localparam VBACK   = 11'd23;
